`timescale 1ns / 1ps

module dadda24x24_sequential(
    input clk,
    input enable,
    input nrst,
    input [23:0] a,
    input [23:0] b,
    output reg [47:0] z,
    output busy,
    output done
    );

    //partial product generator
    parameter N = 24;

    wire ps [N-1:0][N-1:0];
    reg p [N-1:0][N-1:0];

    genvar i;
    genvar j;

    generate
        for (i = 0; i < N; i = i + 1) begin
            for (j = 0; j < N; j = j + 1) begin
                and and0(ps[j][i], a[i], b[j]);
            end
        end
    endgenerate

    wire s [576:0];
    wire c [576:0];

    reg [8:0] counter;
    reg bsy;

    assign busy = bsy;
    assign done = counter[0];

    reg sr [576:0];
    reg cr [576:0];

    wire [(N*2)-2 : 0] result;

    integer x;
    integer y;
    always @(posedge clk, negedge nrst) begin
        if (!nrst) begin
            counter <= 10'd0;
            bsy <= 1'b0;
        end else begin
            counter <= counter >> 1;
          
            if (enable && !bsy) begin
                bsy <= 1'b1;
                counter[8] <= 1'b1;
                for (x = 0; x < N; x = x + 1) begin
                    for (y = 0; y < N; y = y + 1) begin
                        p[y][x] <= ps[y][x];
                    end 
                end
            end

            for (x = 0; x < N*N; x = x + 1) begin
                sr[x] <= s[x];
                cr[x] <= c[x];
            end

            if (counter[1]) begin
                z[(N*2)-1:1] <= result;
                z[0] <= p[0][0];
                bsy <= 1'b0;
            end
        end
    end
//step 6
    ha a0(p[0][19], p[1][18], s[0], c[0]);
    fa a1(p[0][20], p[1][19], p[2][18], s[1], c[1]);
    ha a2(p[3][17], p[4][16], s[2], c[2]);
    fa a3(p[0][21], p[1][20], p[2][19], s[3], c[3]);
    fa a4(p[3][18], p[4][17], p[5][16], s[4], c[4]);
    ha a5(p[6][15], p[7][14], s[5], c[5]);
    fa a6(p[0][22], p[1][21], p[2][20], s[6], c[6]);
    fa a7(p[3][19], p[4][18], p[5][17], s[7], c[7]);
    fa a8(p[6][16], p[7][15], p[8][14], s[8], c[8]);
    ha a9(p[9][13], p[10][12], s[9], c[9]);
    fa a10(p[0][23], p[1][22], p[2][21], s[10], c[10]);
    fa a11(p[3][20], p[4][19], p[5][18], s[11], c[11]);
    fa a12(p[6][17], p[7][16], p[8][15], s[12], c[12]);
    fa a13(p[9][14], p[10][13], p[11][12], s[13], c[13]);
    ha a14(p[12][11], p[13][10], s[14], c[14]);
    fa a15(p[1][23], p[2][22], p[3][21], s[15], c[15]);
    fa a16(p[4][20], p[5][19], p[6][18], s[16], c[16]);
    fa a17(p[7][17], p[8][16], p[9][15], s[17], c[17]);
    fa a18(p[10][14], p[11][13], p[12][12], s[18], c[18]);
    ha a19(p[13][11], p[14][10], s[19], c[19]);
    fa a20(p[2][23], p[3][22], p[4][21], s[20], c[20]);
    fa a21(p[5][20], p[6][19], p[7][18], s[21], c[21]);
    fa a22(p[8][17], p[9][16], p[10][15], s[22], c[22]);
    fa a23(p[11][14], p[12][13], p[13][12], s[23], c[23]);
    fa a24(p[3][23], p[4][22], p[5][21], s[24], c[24]);
    fa a25(p[6][20], p[7][19], p[8][18], s[25], c[25]);
    fa a26(p[9][17], p[10][16], p[11][15], s[26], c[26]);
    fa a27(p[4][23], p[5][22], p[6][21], s[27], c[27]);
    fa a28(p[7][20], p[8][19], p[9][18], s[28], c[28]);
    fa a29(p[5][23], p[6][22], p[7][21], s[29], c[29]);
//step 5
    ha a30(p[0][13], p[1][12], s[30], c[30]);
    fa a31(p[0][14], p[1][13], p[2][12], s[31], c[31]);
    ha a32(p[3][11], p[4][10], s[32], c[32]);
    fa a33(p[0][15], p[1][14], p[2][13], s[33], c[33]);
    fa a34(p[3][12], p[4][11], p[5][10], s[34], c[34]);
    ha a35(p[6][9], p[7][8], s[35], c[35]);
    fa a36(p[0][16], p[1][15], p[2][14], s[36], c[36]);
    fa a37(p[3][13], p[4][12], p[5][11], s[37], c[37]);
    fa a38(p[6][10], p[7][9], p[8][8], s[38], c[38]);
    ha a39(p[9][7], p[10][6], s[39], c[39]);
    fa a40(p[0][17], p[1][16], p[2][15], s[40], c[40]);
    fa a41(p[3][14], p[4][13], p[5][12], s[41], c[41]);
    fa a42(p[6][11], p[7][10], p[8][9], s[42], c[42]);
    fa a43(p[9][8], p[10][7], p[11][6], s[43], c[43]);
    ha a44(p[12][5], p[13][4], s[44], c[44]);
    fa a45(p[0][18], p[1][17], p[2][16], s[45], c[45]);
    fa a46(p[3][15], p[4][14], p[5][13], s[46], c[46]);
    fa a47(p[6][12], p[7][11], p[8][10], s[47], c[47]);
    fa a48(p[9][9], p[10][8], p[11][7], s[48], c[48]);
    fa a49(p[12][6], p[13][5], p[14][4], s[49], c[49]);
    ha a50(p[15][3], p[16][2], s[50], c[50]);
    fa a51(p[2][17], p[3][16], p[4][15], s[51], c[51]);
    fa a52(p[5][14], p[6][13], p[7][12], s[52], c[52]);
    fa a53(p[8][11], p[9][10], p[10][9], s[53], c[53]);
    fa a54(p[11][8], p[12][7], p[13][6], s[54], c[54]);
    fa a55(p[14][5], p[15][4], p[16][3], s[55], c[55]);
    fa a56(p[17][2], p[18][1], p[19][0], s[56], c[56]);
    fa a57(p[5][15], p[6][14], p[7][13], s[57], c[57]);
    fa a58(p[8][12], p[9][11], p[10][10], s[58], c[58]);
    fa a59(p[11][9], p[12][8], p[13][7], s[59], c[59]);
    fa a60(p[14][6], p[15][5], p[16][4], s[60], c[60]);
    fa a61(p[17][3], p[18][2], p[19][1], s[61], c[61]);
    fa a62(p[20][0], cr[0], sr[1], s[62], c[62]);
    fa a63(p[8][13], p[9][12], p[10][11], s[63], c[63]);
    fa a64(p[11][10], p[12][9], p[13][8], s[64], c[64]);
    fa a65(p[14][7], p[15][6], p[16][5], s[65], c[65]);
    fa a66(p[17][4], p[18][3], p[19][2], s[66], c[66]);
    fa a67(p[20][1], p[21][0], cr[1], s[67], c[67]);
    fa a68(cr[2], sr[3], sr[4], s[68], c[68]);
    fa a69(p[11][11], p[12][10], p[13][9], s[69], c[69]);
    fa a70(p[14][8], p[15][7], p[16][6], s[70], c[70]);
    fa a71(p[17][5], p[18][4], p[19][3], s[71], c[71]);
    fa a72(p[20][2], p[21][1], p[22][0], s[72], c[72]);
    fa a73(cr[3], cr[4], cr[5], s[73], c[73]);
    fa a74(sr[6], sr[7], sr[8], s[74], c[74]);
    fa a75(p[14][9], p[15][8], p[16][7], s[75], c[75]);
    fa a76(p[17][6], p[18][5], p[19][4], s[76], c[76]);
    fa a77(p[20][3], p[21][2], p[22][1], s[77], c[77]);
    fa a78(p[23][0], cr[6], cr[7], s[78], c[78]);
    fa a79(cr[8], cr[9], sr[10], s[79], c[79]);
    fa a80(sr[11], sr[12], sr[13], s[80], c[80]);
    fa a81(p[15][9], p[16][8], p[17][7], s[81], c[81]);
    fa a82(p[18][6], p[19][5], p[20][4], s[82], c[82]);
    fa a83(p[21][3], p[22][2], p[23][1], s[83], c[83]);
    fa a84(cr[10], cr[11], cr[12], s[84], c[84]);
    fa a85(cr[13], cr[14], sr[15], s[85], c[85]);
    fa a86(sr[16], sr[17], sr[18], s[86], c[86]);
    fa a87(p[14][11], p[15][10], p[16][9], s[87], c[87]);
    fa a88(p[17][8], p[18][7], p[19][6], s[88], c[88]);
    fa a89(p[20][5], p[21][4], p[22][3], s[89], c[89]);
    fa a90(p[23][2], cr[15], cr[16], s[90], c[90]);
    fa a91(cr[17], cr[18], cr[19], s[91], c[91]);
    fa a92(sr[20], sr[21], sr[22], s[92], c[92]);
    fa a93(p[12][14], p[13][13], p[14][12], s[93], c[93]);
    fa a94(p[15][11], p[16][10], p[17][9], s[94], c[94]);
    fa a95(p[18][8], p[19][7], p[20][6], s[95], c[95]);
    fa a96(p[21][5], p[22][4], p[23][3], s[96], c[96]);
    fa a97(cr[20], cr[21], cr[22], s[97], c[97]);
    fa a98(cr[23], sr[24], sr[25], s[98], c[98]);
    fa a99(p[10][17], p[11][16], p[12][15], s[99], c[99]);
    fa a100(p[13][14], p[14][13], p[15][12], s[100], c[100]);
    fa a101(p[16][11], p[17][10], p[18][9], s[101], c[101]);
    fa a102(p[19][8], p[20][7], p[21][6], s[102], c[102]);
    fa a103(p[22][5], p[23][4], cr[24], s[103], c[103]);
    fa a104(cr[25], cr[26], sr[27], s[104], c[104]);
    fa a105(p[8][20], p[9][19], p[10][18], s[105], c[105]);
    fa a106(p[11][17], p[12][16], p[13][15], s[106], c[106]);
    fa a107(p[14][14], p[15][13], p[16][12], s[107], c[107]);
    fa a108(p[17][11], p[18][10], p[19][9], s[108], c[108]);
    fa a109(p[20][8], p[21][7], p[22][6], s[109], c[109]);
    fa a110(p[23][5], cr[27], cr[28], s[110], c[110]);
    fa a111(p[6][23], p[7][22], p[8][21], s[111], c[111]);
    fa a112(p[9][20], p[10][19], p[11][18], s[112], c[112]);
    fa a113(p[12][17], p[13][16], p[14][15], s[113], c[113]);
    fa a114(p[15][14], p[16][13], p[17][12], s[114], c[114]);
    fa a115(p[18][11], p[19][10], p[20][9], s[115], c[115]);
    fa a116(p[21][8], p[22][7], p[23][6], s[116], c[116]);
    fa a117(p[7][23], p[8][22], p[9][21], s[117], c[117]);
    fa a118(p[10][20], p[11][19], p[12][18], s[118], c[118]);
    fa a119(p[13][17], p[14][16], p[15][15], s[119], c[119]);
    fa a120(p[16][14], p[17][13], p[18][12], s[120], c[120]);
    fa a121(p[19][11], p[20][10], p[21][9], s[121], c[121]);
    fa a122(p[8][23], p[9][22], p[10][21], s[122], c[122]);
    fa a123(p[11][20], p[12][19], p[13][18], s[123], c[123]);
    fa a124(p[14][17], p[15][16], p[16][15], s[124], c[124]);
    fa a125(p[17][14], p[18][13], p[19][12], s[125], c[125]);
    fa a126(p[9][23], p[10][22], p[11][21], s[126], c[126]);
    fa a127(p[12][20], p[13][19], p[14][18], s[127], c[127]);
    fa a128(p[15][17], p[16][16], p[17][15], s[128], c[128]);
    fa a129(p[10][23], p[11][22], p[12][21], s[129], c[129]);
    fa a130(p[13][20], p[14][19], p[15][18], s[130], c[130]);
    fa a131(p[11][23], p[12][22], p[13][21], s[131], c[131]);
//step 4
    ha a132(p[0][9], p[1][8], s[132], c[132]);
    fa a133(p[0][10], p[1][9], p[2][8], s[133], c[133]);
    ha a134(p[3][7], p[4][6], s[134], c[134]);
    fa a135(p[0][11], p[1][10], p[2][9], s[135], c[135]);
    fa a136(p[3][8], p[4][7], p[5][6], s[136], c[136]);
    ha a137(p[6][5], p[7][4], s[137], c[137]);
    fa a138(p[0][12], p[1][11], p[2][10], s[138], c[138]);
    fa a139(p[3][9], p[4][8], p[5][7], s[139], c[139]);
    fa a140(p[6][6], p[7][5], p[8][4], s[140], c[140]);
    ha a141(p[9][3], p[10][2], s[141], c[141]);
    fa a142(p[2][11], p[3][10], p[4][9], s[142], c[142]);
    fa a143(p[5][8], p[6][7], p[7][6], s[143], c[143]);
    fa a144(p[8][5], p[9][4], p[10][3], s[144], c[144]);
    fa a145(p[11][2], p[12][1], p[13][0], s[145], c[145]);
    fa a146(p[5][9], p[6][8], p[7][7], s[146], c[146]);
    fa a147(p[8][6], p[9][5], p[10][4], s[147], c[147]);
    fa a148(p[11][3], p[12][2], p[13][1], s[148], c[148]);
    fa a149(p[14][0], cr[30], sr[31], s[149], c[149]);
    fa a150(p[8][7], p[9][6], p[10][5], s[150], c[150]);
    fa a151(p[11][4], p[12][3], p[13][2], s[151], c[151]);
    fa a152(p[14][1], p[15][0], cr[31], s[152], c[152]);
    fa a153(cr[32], sr[33], sr[34], s[153], c[153]);
    fa a154(p[11][5], p[12][4], p[13][3], s[154], c[154]);
    fa a155(p[14][2], p[15][1], p[16][0], s[155], c[155]);
    fa a156(cr[33], cr[34], cr[35], s[156], c[156]);
    fa a157(sr[36], sr[37], sr[38], s[157], c[157]);
    fa a158(p[14][3], p[15][2], p[16][1], s[158], c[158]);
    fa a159(p[17][0], cr[36], cr[37], s[159], c[159]);
    fa a160(cr[38], cr[39], sr[40], s[160], c[160]);
    fa a161(sr[41], sr[42], sr[43], s[161], c[161]);
    fa a162(p[17][1], p[18][0], cr[40], s[162], c[162]);
    fa a163(cr[41], cr[42], cr[43], s[163], c[163]);
    fa a164(cr[44], sr[45], sr[46], s[164], c[164]);
    fa a165(sr[47], sr[48], sr[49], s[165], c[165]);
    fa a166(sr[0], cr[45], cr[46], s[166], c[166]);
    fa a167(cr[47], cr[48], cr[49], s[167], c[167]);
    fa a168(cr[50], sr[51], sr[52], s[168], c[168]);
    fa a169(sr[53], sr[54], sr[55], s[169], c[169]);
    fa a170(sr[2], cr[51], cr[52], s[170], c[170]);
    fa a171(cr[53], cr[54], cr[55], s[171], c[171]);
    fa a172(cr[56], sr[57], sr[58], s[172], c[172]);
    fa a173(sr[59], sr[60], sr[61], s[173], c[173]);
    fa a174(sr[5], cr[57], cr[58], s[174], c[174]);
    fa a175(cr[59], cr[60], cr[61], s[175], c[175]);
    fa a176(cr[62], sr[63], sr[64], s[176], c[176]);
    fa a177(sr[65], sr[66], sr[67], s[177], c[177]);
    fa a178(sr[9], cr[63], cr[64], s[178], c[178]);
    fa a179(cr[65], cr[66], cr[67], s[179], c[179]);
    fa a180(cr[68], sr[69], sr[70], s[180], c[180]);
    fa a181(sr[71], sr[72], sr[73], s[181], c[181]);
    fa a182(sr[14], cr[69], cr[70], s[182], c[182]);
    fa a183(cr[71], cr[72], cr[73], s[183], c[183]);
    fa a184(cr[74], sr[75], sr[76], s[184], c[184]);
    fa a185(sr[77], sr[78], sr[79], s[185], c[185]);
    fa a186(sr[19], cr[75], cr[76], s[186], c[186]);
    fa a187(cr[77], cr[78], cr[79], s[187], c[187]);
    fa a188(cr[80], sr[81], sr[82], s[188], c[188]);
    fa a189(sr[83], sr[84], sr[85], s[189], c[189]);
    fa a190(sr[23], cr[81], cr[82], s[190], c[190]);
    fa a191(cr[83], cr[84], cr[85], s[191], c[191]);
    fa a192(cr[86], sr[87], sr[88], s[192], c[192]);
    fa a193(sr[89], sr[90], sr[91], s[193], c[193]);
    fa a194(sr[26], cr[87], cr[88], s[194], c[194]);
    fa a195(cr[89], cr[90], cr[91], s[195], c[195]);
    fa a196(cr[92], sr[93], sr[94], s[196], c[196]);
    fa a197(sr[95], sr[96], sr[97], s[197], c[197]);
    fa a198(sr[28], cr[93], cr[94], s[198], c[198]);
    fa a199(cr[95], cr[96], cr[97], s[199], c[199]);
    fa a200(cr[98], sr[99], sr[100], s[200], c[200]);
    fa a201(sr[101], sr[102], sr[103], s[201], c[201]);
    fa a202(sr[29], cr[99], cr[100], s[202], c[202]);
    fa a203(cr[101], cr[102], cr[103], s[203], c[203]);
    fa a204(cr[104], sr[105], sr[106], s[204], c[204]);
    fa a205(sr[107], sr[108], sr[109], s[205], c[205]);
    fa a206(cr[29], cr[105], cr[106], s[206], c[206]);
    fa a207(cr[107], cr[108], cr[109], s[207], c[207]);
    fa a208(cr[110], sr[111], sr[112], s[208], c[208]);
    fa a209(sr[113], sr[114], sr[115], s[209], c[209]);
    fa a210(p[22][8], p[23][7], cr[111], s[210], c[210]);
    fa a211(cr[112], cr[113], cr[114], s[211], c[211]);
    fa a212(cr[115], cr[116], sr[117], s[212], c[212]);
    fa a213(sr[118], sr[119], sr[120], s[213], c[213]);
    fa a214(p[20][11], p[21][10], p[22][9], s[214], c[214]);
    fa a215(p[23][8], cr[117], cr[118], s[215], c[215]);
    fa a216(cr[119], cr[120], cr[121], s[216], c[216]);
    fa a217(sr[122], sr[123], sr[124], s[217], c[217]);
    fa a218(p[18][14], p[19][13], p[20][12], s[218], c[218]);
    fa a219(p[21][11], p[22][10], p[23][9], s[219], c[219]);
    fa a220(cr[122], cr[123], cr[124], s[220], c[220]);
    fa a221(cr[125], sr[126], sr[127], s[221], c[221]);
    fa a222(p[16][17], p[17][16], p[18][15], s[222], c[222]);
    fa a223(p[19][14], p[20][13], p[21][12], s[223], c[223]);
    fa a224(p[22][11], p[23][10], cr[126], s[224], c[224]);
    fa a225(cr[127], cr[128], sr[129], s[225], c[225]);
    fa a226(p[14][20], p[15][19], p[16][18], s[226], c[226]);
    fa a227(p[17][17], p[18][16], p[19][15], s[227], c[227]);
    fa a228(p[20][14], p[21][13], p[22][12], s[228], c[228]);
    fa a229(p[23][11], cr[129], cr[130], s[229], c[229]);
    fa a230(p[12][23], p[13][22], p[14][21], s[230], c[230]);
    fa a231(p[15][20], p[16][19], p[17][18], s[231], c[231]);
    fa a232(p[18][17], p[19][16], p[20][15], s[232], c[232]);
    fa a233(p[21][14], p[22][13], p[23][12], s[233], c[233]);
    fa a234(p[13][23], p[14][22], p[15][21], s[234], c[234]);
    fa a235(p[16][20], p[17][19], p[18][18], s[235], c[235]);
    fa a236(p[19][17], p[20][16], p[21][15], s[236], c[236]);
    fa a237(p[14][23], p[15][22], p[16][21], s[237], c[237]);
    fa a238(p[17][20], p[18][19], p[19][18], s[238], c[238]);
    fa a239(p[15][23], p[16][22], p[17][21], s[239], c[239]);
//step 3
    ha a240(p[0][6], p[1][5], s[240], c[240]);
    fa a241(p[0][7], p[1][6], p[2][5], s[241], c[241]);
    ha a242(p[3][4], p[4][3], s[242], c[242]);
    fa a243(p[0][8], p[1][7], p[2][6], s[243], c[243]);
    fa a244(p[3][5], p[4][4], p[5][3], s[244], c[244]);
    ha a245(p[6][2], p[7][1], s[245], c[245]);
    fa a246(p[2][7], p[3][6], p[4][5], s[246], c[246]);
    fa a247(p[5][4], p[6][3], p[7][2], s[247], c[247]);
    fa a248(p[8][1], p[9][0], sr[132], s[248], c[248]);
    fa a249(p[5][5], p[6][4], p[7][3], s[249], c[249]);
    fa a250(p[8][2], p[9][1], p[10][0], s[250], c[250]);
    fa a251(cr[132], sr[133], sr[134], s[251], c[251]);
    fa a252(p[8][3], p[9][2], p[10][1], s[252], c[252]);
    fa a253(p[11][0], cr[133], cr[134], s[253], c[253]);
    fa a254(sr[135], sr[136], sr[137], s[254], c[254]);
    fa a255(p[11][1], p[12][0], cr[135], s[255], c[255]);
    fa a256(cr[136], cr[137], sr[138], s[256], c[256]);
    fa a257(sr[139], sr[140], sr[141], s[257], c[257]);
    fa a258(sr[30], cr[138], cr[139], s[258], c[258]);
    fa a259(cr[140], cr[141], sr[142], s[259], c[259]);
    fa a260(sr[143], sr[144], sr[145], s[260], c[260]);
    fa a261(sr[32], cr[142], cr[143], s[261], c[261]);
    fa a262(cr[144], cr[145], sr[146], s[262], c[262]);
    fa a263(sr[147], sr[148], sr[149], s[263], c[263]);
    fa a264(sr[35], cr[146], cr[147], s[264], c[264]);
    fa a265(cr[148], cr[149], sr[150], s[265], c[265]);
    fa a266(sr[151], sr[152], sr[153], s[266], c[266]);
    fa a267(sr[39], cr[150], cr[151], s[267], c[267]);
    fa a268(cr[152], cr[153], sr[154], s[268], c[268]);
    fa a269(sr[155], sr[156], sr[157], s[269], c[269]);
    fa a270(sr[44], cr[154], cr[155], s[270], c[270]);
    fa a271(cr[156], cr[157], sr[158], s[271], c[271]);
    fa a272(sr[159], sr[160], sr[161], s[272], c[272]);
    fa a273(sr[50], cr[158], cr[159], s[273], c[273]);
    fa a274(cr[160], cr[161], sr[162], s[274], c[274]);
    fa a275(sr[163], sr[164], sr[165], s[275], c[275]);
    fa a276(sr[56], cr[162], cr[163], s[276], c[276]);
    fa a277(cr[164], cr[165], sr[166], s[277], c[277]);
    fa a278(sr[167], sr[168], sr[169], s[278], c[278]);
    fa a279(sr[62], cr[166], cr[167], s[279], c[279]);
    fa a280(cr[168], cr[169], sr[170], s[280], c[280]);
    fa a281(sr[171], sr[172], sr[173], s[281], c[281]);
    fa a282(sr[68], cr[170], cr[171], s[282], c[282]);
    fa a283(cr[172], cr[173], sr[174], s[283], c[283]);
    fa a284(sr[175], sr[176], sr[177], s[284], c[284]);
    fa a285(sr[74], cr[174], cr[175], s[285], c[285]);
    fa a286(cr[176], cr[177], sr[178], s[286], c[286]);
    fa a287(sr[179], sr[180], sr[181], s[287], c[287]);
    fa a288(sr[80], cr[178], cr[179], s[288], c[288]);
    fa a289(cr[180], cr[181], sr[182], s[289], c[289]);
    fa a290(sr[183], sr[184], sr[185], s[290], c[290]);
    fa a291(sr[86], cr[182], cr[183], s[291], c[291]);
    fa a292(cr[184], cr[185], sr[186], s[292], c[292]);
    fa a293(sr[187], sr[188], sr[189], s[293], c[293]);
    fa a294(sr[92], cr[186], cr[187], s[294], c[294]);
    fa a295(cr[188], cr[189], sr[190], s[295], c[295]);
    fa a296(sr[191], sr[192], sr[193], s[296], c[296]);
    fa a297(sr[98], cr[190], cr[191], s[297], c[297]);
    fa a298(cr[192], cr[193], sr[194], s[298], c[298]);
    fa a299(sr[195], sr[196], sr[197], s[299], c[299]);
    fa a300(sr[104], cr[194], cr[195], s[300], c[300]);
    fa a301(cr[196], cr[197], sr[198], s[301], c[301]);
    fa a302(sr[199], sr[200], sr[201], s[302], c[302]);
    fa a303(sr[110], cr[198], cr[199], s[303], c[303]);
    fa a304(cr[200], cr[201], sr[202], s[304], c[304]);
    fa a305(sr[203], sr[204], sr[205], s[305], c[305]);
    fa a306(sr[116], cr[202], cr[203], s[306], c[306]);
    fa a307(cr[204], cr[205], sr[206], s[307], c[307]);
    fa a308(sr[207], sr[208], sr[209], s[308], c[308]);
    fa a309(sr[121], cr[206], cr[207], s[309], c[309]);
    fa a310(cr[208], cr[209], sr[210], s[310], c[310]);
    fa a311(sr[211], sr[212], sr[213], s[311], c[311]);
    fa a312(sr[125], cr[210], cr[211], s[312], c[312]);
    fa a313(cr[212], cr[213], sr[214], s[313], c[313]);
    fa a314(sr[215], sr[216], sr[217], s[314], c[314]);
    fa a315(sr[128], cr[214], cr[215], s[315], c[315]);
    fa a316(cr[216], cr[217], sr[218], s[316], c[316]);
    fa a317(sr[219], sr[220], sr[221], s[317], c[317]);
    fa a318(sr[130], cr[218], cr[219], s[318], c[318]);
    fa a319(cr[220], cr[221], sr[222], s[319], c[319]);
    fa a320(sr[223], sr[224], sr[225], s[320], c[320]);
    fa a321(sr[131], cr[222], cr[223], s[321], c[321]);
    fa a322(cr[224], cr[225], sr[226], s[322], c[322]);
    fa a323(sr[227], sr[228], sr[229], s[323], c[323]);
    fa a324(cr[131], cr[226], cr[227], s[324], c[324]);
    fa a325(cr[228], cr[229], sr[230], s[325], c[325]);
    fa a326(sr[231], sr[232], sr[233], s[326], c[326]);
    fa a327(p[22][14], p[23][13], cr[230], s[327], c[327]);
    fa a328(cr[231], cr[232], cr[233], s[328], c[328]);
    fa a329(sr[234], sr[235], sr[236], s[329], c[329]);
    fa a330(p[20][17], p[21][16], p[22][15], s[330], c[330]);
    fa a331(p[23][14], cr[234], cr[235], s[331], c[331]);
    fa a332(cr[236], sr[237], sr[238], s[332], c[332]);
    fa a333(p[18][20], p[19][19], p[20][18], s[333], c[333]);
    fa a334(p[21][17], p[22][16], p[23][15], s[334], c[334]);
    fa a335(cr[237], cr[238], sr[239], s[335], c[335]);
    fa a336(p[16][23], p[17][22], p[18][21], s[336], c[336]);
    fa a337(p[19][20], p[20][19], p[21][18], s[337], c[337]);
    fa a338(p[22][17], p[23][16], cr[239], s[338], c[338]);
    fa a339(p[17][23], p[18][22], p[19][21], s[339], c[339]);
    fa a340(p[20][20], p[21][19], p[22][18], s[340], c[340]);
    fa a341(p[18][23], p[19][22], p[20][21], s[341], c[341]);
//step 2
    ha a342(p[0][4], p[1][3], s[342], c[342]);
    fa a343(p[0][5], p[1][4], p[2][3], s[343], c[343]);
    ha a344(p[3][2], p[4][1], s[344], c[344]);
    fa a345(p[2][4], p[3][3], p[4][2], s[345], c[345]);
    fa a346(p[5][1], p[6][0], sr[240], s[346], c[346]);
    fa a347(p[5][2], p[6][1], p[7][0], s[347], c[347]);
    fa a348(cr[240], sr[241], sr[242], s[348], c[348]);
    fa a349(p[8][0], cr[241], cr[242], s[349], c[349]);
    fa a350(sr[243], sr[244], sr[245], s[350], c[350]);
    fa a351(cr[243], cr[244], cr[245], s[351], c[351]);
    fa a352(sr[246], sr[247], sr[248], s[352], c[352]);
    fa a353(cr[246], cr[247], cr[248], s[353], c[353]);
    fa a354(sr[249], sr[250], sr[251], s[354], c[354]);
    fa a355(cr[249], cr[250], cr[251], s[355], c[355]);
    fa a356(sr[252], sr[253], sr[254], s[356], c[356]);
    fa a357(cr[252], cr[253], cr[254], s[357], c[357]);
    fa a358(sr[255], sr[256], sr[257], s[358], c[358]);
    fa a359(cr[255], cr[256], cr[257], s[359], c[359]);
    fa a360(sr[258], sr[259], sr[260], s[360], c[360]);
    fa a361(cr[258], cr[259], cr[260], s[361], c[361]);
    fa a362(sr[261], sr[262], sr[263], s[362], c[362]);
    fa a363(cr[261], cr[262], cr[263], s[363], c[363]);
    fa a364(sr[264], sr[265], sr[266], s[364], c[364]);
    fa a365(cr[264], cr[265], cr[266], s[365], c[365]);
    fa a366(sr[267], sr[268], sr[269], s[366], c[366]);
    fa a367(cr[267], cr[268], cr[269], s[367], c[367]);
    fa a368(sr[270], sr[271], sr[272], s[368], c[368]);
    fa a369(cr[270], cr[271], cr[272], s[369], c[369]);
    fa a370(sr[273], sr[274], sr[275], s[370], c[370]);
    fa a371(cr[273], cr[274], cr[275], s[371], c[371]);
    fa a372(sr[276], sr[277], sr[278], s[372], c[372]);
    fa a373(cr[276], cr[277], cr[278], s[373], c[373]);
    fa a374(sr[279], sr[280], sr[281], s[374], c[374]);
    fa a375(cr[279], cr[280], cr[281], s[375], c[375]);
    fa a376(sr[282], sr[283], sr[284], s[376], c[376]);
    fa a377(cr[282], cr[283], cr[284], s[377], c[377]);
    fa a378(sr[285], sr[286], sr[287], s[378], c[378]);
    fa a379(cr[285], cr[286], cr[287], s[379], c[379]);
    fa a380(sr[288], sr[289], sr[290], s[380], c[380]);
    fa a381(cr[288], cr[289], cr[290], s[381], c[381]);
    fa a382(sr[291], sr[292], sr[293], s[382], c[382]);
    fa a383(cr[291], cr[292], cr[293], s[383], c[383]);
    fa a384(sr[294], sr[295], sr[296], s[384], c[384]);
    fa a385(cr[294], cr[295], cr[296], s[385], c[385]);
    fa a386(sr[297], sr[298], sr[299], s[386], c[386]);
    fa a387(cr[297], cr[298], cr[299], s[387], c[387]);
    fa a388(sr[300], sr[301], sr[302], s[388], c[388]);
    fa a389(cr[300], cr[301], cr[302], s[389], c[389]);
    fa a390(sr[303], sr[304], sr[305], s[390], c[390]);
    fa a391(cr[303], cr[304], cr[305], s[391], c[391]);
    fa a392(sr[306], sr[307], sr[308], s[392], c[392]);
    fa a393(cr[306], cr[307], cr[308], s[393], c[393]);
    fa a394(sr[309], sr[310], sr[311], s[394], c[394]);
    fa a395(cr[309], cr[310], cr[311], s[395], c[395]);
    fa a396(sr[312], sr[313], sr[314], s[396], c[396]);
    fa a397(cr[312], cr[313], cr[314], s[397], c[397]);
    fa a398(sr[315], sr[316], sr[317], s[398], c[398]);
    fa a399(cr[315], cr[316], cr[317], s[399], c[399]);
    fa a400(sr[318], sr[319], sr[320], s[400], c[400]);
    fa a401(cr[318], cr[319], cr[320], s[401], c[401]);
    fa a402(sr[321], sr[322], sr[323], s[402], c[402]);
    fa a403(cr[321], cr[322], cr[323], s[403], c[403]);
    fa a404(sr[324], sr[325], sr[326], s[404], c[404]);
    fa a405(cr[324], cr[325], cr[326], s[405], c[405]);
    fa a406(sr[327], sr[328], sr[329], s[406], c[406]);
    fa a407(cr[327], cr[328], cr[329], s[407], c[407]);
    fa a408(sr[330], sr[331], sr[332], s[408], c[408]);
    fa a409(cr[330], cr[331], cr[332], s[409], c[409]);
    fa a410(sr[333], sr[334], sr[335], s[410], c[410]);
    fa a411(cr[333], cr[334], cr[335], s[411], c[411]);
    fa a412(sr[336], sr[337], sr[338], s[412], c[412]);
    fa a413(p[23][17], cr[336], cr[337], s[413], c[413]);
    fa a414(cr[338], sr[339], sr[340], s[414], c[414]);
    fa a415(p[21][20], p[22][19], p[23][18], s[415], c[415]);
    fa a416(cr[339], cr[340], sr[341], s[416], c[416]);
    fa a417(p[19][23], p[20][22], p[21][21], s[417], c[417]);
    fa a418(p[22][20], p[23][19], cr[341], s[418], c[418]);
    fa a419(p[20][23], p[21][22], p[22][21], s[419], c[419]);
//step 1
    ha a420(p[0][3], p[1][2], s[420], c[420]);
    fa a421(p[2][2], p[3][1], p[4][0], s[421], c[421]);
    fa a422(p[5][0], cr[342], sr[343], s[422], c[422]);
    fa a423(cr[343], cr[344], sr[345], s[423], c[423]);
    fa a424(cr[345], cr[346], sr[347], s[424], c[424]);
    fa a425(cr[347], cr[348], sr[349], s[425], c[425]);
    fa a426(cr[349], cr[350], sr[351], s[426], c[426]);
    fa a427(cr[351], cr[352], sr[353], s[427], c[427]);
    fa a428(cr[353], cr[354], sr[355], s[428], c[428]);
    fa a429(cr[355], cr[356], sr[357], s[429], c[429]);
    fa a430(cr[357], cr[358], sr[359], s[430], c[430]);
    fa a431(cr[359], cr[360], sr[361], s[431], c[431]);
    fa a432(cr[361], cr[362], sr[363], s[432], c[432]);
    fa a433(cr[363], cr[364], sr[365], s[433], c[433]);
    fa a434(cr[365], cr[366], sr[367], s[434], c[434]);
    fa a435(cr[367], cr[368], sr[369], s[435], c[435]);
    fa a436(cr[369], cr[370], sr[371], s[436], c[436]);
    fa a437(cr[371], cr[372], sr[373], s[437], c[437]);
    fa a438(cr[373], cr[374], sr[375], s[438], c[438]);
    fa a439(cr[375], cr[376], sr[377], s[439], c[439]);
    fa a440(cr[377], cr[378], sr[379], s[440], c[440]);
    fa a441(cr[379], cr[380], sr[381], s[441], c[441]);
    fa a442(cr[381], cr[382], sr[383], s[442], c[442]);
    fa a443(cr[383], cr[384], sr[385], s[443], c[443]);
    fa a444(cr[385], cr[386], sr[387], s[444], c[444]);
    fa a445(cr[387], cr[388], sr[389], s[445], c[445]);
    fa a446(cr[389], cr[390], sr[391], s[446], c[446]);
    fa a447(cr[391], cr[392], sr[393], s[447], c[447]);
    fa a448(cr[393], cr[394], sr[395], s[448], c[448]);
    fa a449(cr[395], cr[396], sr[397], s[449], c[449]);
    fa a450(cr[397], cr[398], sr[399], s[450], c[450]);
    fa a451(cr[399], cr[400], sr[401], s[451], c[451]);
    fa a452(cr[401], cr[402], sr[403], s[452], c[452]);
    fa a453(cr[403], cr[404], sr[405], s[453], c[453]);
    fa a454(cr[405], cr[406], sr[407], s[454], c[454]);
    fa a455(cr[407], cr[408], sr[409], s[455], c[455]);
    fa a456(cr[409], cr[410], sr[411], s[456], c[456]);
    fa a457(cr[411], cr[412], sr[413], s[457], c[457]);
    fa a458(cr[413], cr[414], sr[415], s[458], c[458]);
    fa a459(cr[415], cr[416], sr[417], s[459], c[459]);
    fa a460(p[23][20], cr[417], cr[418], s[460], c[460]);
    fa a461(p[21][23], p[22][22], p[23][21], s[461], c[461]);
//step 0
    ha a462(p[0][2], p[1][1], s[462], c[462]);
    fa a463(p[2][1], p[3][0], sr[420], s[463], c[463]);
    fa a464(sr[342], cr[420], sr[421], s[464], c[464]);
    fa a465(sr[344], cr[421], sr[422], s[465], c[465]);
    fa a466(sr[346], cr[422], sr[423], s[466], c[466]);
    fa a467(sr[348], cr[423], sr[424], s[467], c[467]);
    fa a468(sr[350], cr[424], sr[425], s[468], c[468]);
    fa a469(sr[352], cr[425], sr[426], s[469], c[469]);
    fa a470(sr[354], cr[426], sr[427], s[470], c[470]);
    fa a471(sr[356], cr[427], sr[428], s[471], c[471]);
    fa a472(sr[358], cr[428], sr[429], s[472], c[472]);
    fa a473(sr[360], cr[429], sr[430], s[473], c[473]);
    fa a474(sr[362], cr[430], sr[431], s[474], c[474]);
    fa a475(sr[364], cr[431], sr[432], s[475], c[475]);
    fa a476(sr[366], cr[432], sr[433], s[476], c[476]);
    fa a477(sr[368], cr[433], sr[434], s[477], c[477]);
    fa a478(sr[370], cr[434], sr[435], s[478], c[478]);
    fa a479(sr[372], cr[435], sr[436], s[479], c[479]);
    fa a480(sr[374], cr[436], sr[437], s[480], c[480]);
    fa a481(sr[376], cr[437], sr[438], s[481], c[481]);
    fa a482(sr[378], cr[438], sr[439], s[482], c[482]);
    fa a483(sr[380], cr[439], sr[440], s[483], c[483]);
    fa a484(sr[382], cr[440], sr[441], s[484], c[484]);
    fa a485(sr[384], cr[441], sr[442], s[485], c[485]);
    fa a486(sr[386], cr[442], sr[443], s[486], c[486]);
    fa a487(sr[388], cr[443], sr[444], s[487], c[487]);
    fa a488(sr[390], cr[444], sr[445], s[488], c[488]);
    fa a489(sr[392], cr[445], sr[446], s[489], c[489]);
    fa a490(sr[394], cr[446], sr[447], s[490], c[490]);
    fa a491(sr[396], cr[447], sr[448], s[491], c[491]);
    fa a492(sr[398], cr[448], sr[449], s[492], c[492]);
    fa a493(sr[400], cr[449], sr[450], s[493], c[493]);
    fa a494(sr[402], cr[450], sr[451], s[494], c[494]);
    fa a495(sr[404], cr[451], sr[452], s[495], c[495]);
    fa a496(sr[406], cr[452], sr[453], s[496], c[496]);
    fa a497(sr[408], cr[453], sr[454], s[497], c[497]);
    fa a498(sr[410], cr[454], sr[455], s[498], c[498]);
    fa a499(sr[412], cr[455], sr[456], s[499], c[499]);
    fa a500(sr[414], cr[456], sr[457], s[500], c[500]);
    fa a501(sr[416], cr[457], sr[458], s[501], c[501]);
    fa a502(sr[418], cr[458], sr[459], s[502], c[502]);
    fa a503(sr[419], cr[459], sr[460], s[503], c[503]);
    fa a504(cr[419], cr[460], sr[461], s[504], c[504]);
    fa a505(p[22][23], p[23][22], cr[461], s[505], c[505]);

    wire[(N*2)-3 : 0] n1;
    wire[(N*2)-3 : 0] n2;
    assign n1[0] = p[0][1];
    assign n1[1] = p[2][0];
    assign n1[2] = cr[462];
    assign n1[3] = cr[463];
    assign n1[4] = cr[464];
    assign n1[5] = cr[465];
    assign n1[6] = cr[466];
    assign n1[7] = cr[467];
    assign n1[8] = cr[468];
    assign n1[9] = cr[469];
    assign n1[10] = cr[470];
    assign n1[11] = cr[471];
    assign n1[12] = cr[472];
    assign n1[13] = cr[473];
    assign n1[14] = cr[474];
    assign n1[15] = cr[475];
    assign n1[16] = cr[476];
    assign n1[17] = cr[477];
    assign n1[18] = cr[478];
    assign n1[19] = cr[479];
    assign n1[20] = cr[480];
    assign n1[21] = cr[481];
    assign n1[22] = cr[482];
    assign n1[23] = cr[483];
    assign n1[24] = cr[484];
    assign n1[25] = cr[485];
    assign n1[26] = cr[486];
    assign n1[27] = cr[487];
    assign n1[28] = cr[488];
    assign n1[29] = cr[489];
    assign n1[30] = cr[490];
    assign n1[31] = cr[491];
    assign n1[32] = cr[492];
    assign n1[33] = cr[493];
    assign n1[34] = cr[494];
    assign n1[35] = cr[495];
    assign n1[36] = cr[496];
    assign n1[37] = cr[497];
    assign n1[38] = cr[498];
    assign n1[39] = cr[499];
    assign n1[40] = cr[500];
    assign n1[41] = cr[501];
    assign n1[42] = cr[502];
    assign n1[43] = cr[503];
    assign n1[44] = cr[504];
    assign n1[45] = p[23][23];
    assign n2[0] = p[1][0];
    assign n2[1] = sr[462];
    assign n2[2] = sr[463];
    assign n2[3] = sr[464];
    assign n2[4] = sr[465];
    assign n2[5] = sr[466];
    assign n2[6] = sr[467];
    assign n2[7] = sr[468];
    assign n2[8] = sr[469];
    assign n2[9] = sr[470];
    assign n2[10] = sr[471];
    assign n2[11] = sr[472];
    assign n2[12] = sr[473];
    assign n2[13] = sr[474];
    assign n2[14] = sr[475];
    assign n2[15] = sr[476];
    assign n2[16] = sr[477];
    assign n2[17] = sr[478];
    assign n2[18] = sr[479];
    assign n2[19] = sr[480];
    assign n2[20] = sr[481];
    assign n2[21] = sr[482];
    assign n2[22] = sr[483];
    assign n2[23] = sr[484];
    assign n2[24] = sr[485];
    assign n2[25] = sr[486];
    assign n2[26] = sr[487];
    assign n2[27] = sr[488];
    assign n2[28] = sr[489];
    assign n2[29] = sr[490];
    assign n2[30] = sr[491];
    assign n2[31] = sr[492];
    assign n2[32] = sr[493];
    assign n2[33] = sr[494];
    assign n2[34] = sr[495];
    assign n2[35] = sr[496];
    assign n2[36] = sr[497];
    assign n2[37] = sr[498];
    assign n2[38] = sr[499];
    assign n2[39] = sr[500];
    assign n2[40] = sr[501];
    assign n2[41] = sr[502];
    assign n2[42] = sr[503];
    assign n2[43] = sr[504];
    assign n2[44] = sr[505];
    assign n2[45] = cr[505];

    assign result = n1+n2;
endmodule
